/////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Behavioral 16-bits multiplier
/////////////////////////////////////////////////////////////////////////////////////////////////////////////

module multiplier_16x16(a, b, out);
    
    output  [31:0]  out;

    input   [15:0]  a; 
    input   [15:0]  b;

    assign out = a * b;

endmodule