////////////////////////////////////////////////////////////////////////
//	Jul 28 2018
//	Transaction fot seq_adder_tb
//	by VAL
////////////////////////////////////////////////////////////////////////

class transaction;

endclass
