/////////////////////////////////////////////////////////////////////////////////////////////////////////////
//  Interrup controller
//  Interrapt controller for My MIPS32_PPL realization
//
//  Author      : VAL
//  Written     : 24 May 2019
//
/////////////////////////////////////////////////////////////////////////////////////////////////////////////

module interrupt_controller();
  
  
  
  
endmodule