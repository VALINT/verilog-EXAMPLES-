///////////////////////////////////////////////////////////////////////////////////////////////////////////////
// 32-bits acumulator
///////////////////////////////////////////////////////////////////////////////////////////////////////////////

module accumulator(in, out, clk, rstb);

output reg  [31:0]  out;

input   [31:0]  in;
input           clk;
input           rstb;

always @(posedge clk or negedge rstb) 
begin
    if(!rstb)
        out <= 'h00000000;
    else
        out <= in;
end

endmodule