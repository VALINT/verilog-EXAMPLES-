////////////////////////////////////////////////////////////////////////
//	Jul 28 2018
//	Environment fot seq_adder_tb
//	by VAL
////////////////////////////////////////////////////////////////////////

interface intf;
	logic			clk;
	logic			rst
	logic	[7:0]	termA;
	logic	[7:0]	termB;
	logic	[7:0]	sum;
	logic			carry;
endinterface
